../delay/delay_pkg.vhd