../delay/delay.vhd